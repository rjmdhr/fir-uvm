package tb_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "agent_config.svh"
	`include "env_config.svh"
	`include "filt_seq_item.svh"
	`include "filt_seq.svh"
	`include "filt_driver.svh"
	`include "filt_scoreboard.svh"
	`include "filt_monitor.svh"
	`include "filt_agent.svh"
	`include "filt_env.svh"
	`include "filt_test.svh"

endpackage